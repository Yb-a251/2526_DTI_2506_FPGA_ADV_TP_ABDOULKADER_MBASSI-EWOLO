// niosv_reset_controller.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module niosv_reset_controller #(
		parameter NUM_RESET_INPUTS          = 2,
		parameter OUTPUT_RESET_SYNC_EDGES   = "deassert",
		parameter SYNC_DEPTH                = 2,
		parameter RESET_REQUEST_PRESENT     = 0,
		parameter RESET_REQ_WAIT_TIME       = 1,
		parameter MIN_RST_ASSERTION_TIME    = 3,
		parameter RESET_REQ_EARLY_DSRT_TIME = 1,
		parameter USE_RESET_REQUEST_IN0     = 0,
		parameter USE_RESET_REQUEST_IN1     = 0,
		parameter USE_RESET_REQUEST_IN2     = 0,
		parameter USE_RESET_REQUEST_IN3     = 0,
		parameter USE_RESET_REQUEST_IN4     = 0,
		parameter USE_RESET_REQUEST_IN5     = 0,
		parameter USE_RESET_REQUEST_IN6     = 0,
		parameter USE_RESET_REQUEST_IN7     = 0,
		parameter USE_RESET_REQUEST_IN8     = 0,
		parameter USE_RESET_REQUEST_IN9     = 0,
		parameter USE_RESET_REQUEST_IN10    = 0,
		parameter USE_RESET_REQUEST_IN11    = 0,
		parameter USE_RESET_REQUEST_IN12    = 0,
		parameter USE_RESET_REQUEST_IN13    = 0,
		parameter USE_RESET_REQUEST_IN14    = 0,
		parameter USE_RESET_REQUEST_IN15    = 0,
		parameter ADAPT_RESET_REQUEST       = 0
	) (
		input  wire  reset_in0, // reset_in0.reset
		input  wire  reset_in1, // reset_in1.reset
		input  wire  clk,       //       clk.clk
		output wire  reset_out  // reset_out.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (NUM_RESET_INPUTS),
		.OUTPUT_RESET_SYNC_EDGES   (OUTPUT_RESET_SYNC_EDGES),
		.SYNC_DEPTH                (SYNC_DEPTH),
		.RESET_REQUEST_PRESENT     (RESET_REQUEST_PRESENT),
		.RESET_REQ_WAIT_TIME       (RESET_REQ_WAIT_TIME),
		.MIN_RST_ASSERTION_TIME    (MIN_RST_ASSERTION_TIME),
		.RESET_REQ_EARLY_DSRT_TIME (RESET_REQ_EARLY_DSRT_TIME),
		.USE_RESET_REQUEST_IN0     (USE_RESET_REQUEST_IN0),
		.USE_RESET_REQUEST_IN1     (USE_RESET_REQUEST_IN1),
		.USE_RESET_REQUEST_IN2     (USE_RESET_REQUEST_IN2),
		.USE_RESET_REQUEST_IN3     (USE_RESET_REQUEST_IN3),
		.USE_RESET_REQUEST_IN4     (USE_RESET_REQUEST_IN4),
		.USE_RESET_REQUEST_IN5     (USE_RESET_REQUEST_IN5),
		.USE_RESET_REQUEST_IN6     (USE_RESET_REQUEST_IN6),
		.USE_RESET_REQUEST_IN7     (USE_RESET_REQUEST_IN7),
		.USE_RESET_REQUEST_IN8     (USE_RESET_REQUEST_IN8),
		.USE_RESET_REQUEST_IN9     (USE_RESET_REQUEST_IN9),
		.USE_RESET_REQUEST_IN10    (USE_RESET_REQUEST_IN10),
		.USE_RESET_REQUEST_IN11    (USE_RESET_REQUEST_IN11),
		.USE_RESET_REQUEST_IN12    (USE_RESET_REQUEST_IN12),
		.USE_RESET_REQUEST_IN13    (USE_RESET_REQUEST_IN13),
		.USE_RESET_REQUEST_IN14    (USE_RESET_REQUEST_IN14),
		.USE_RESET_REQUEST_IN15    (USE_RESET_REQUEST_IN15),
		.ADAPT_RESET_REQUEST       (ADAPT_RESET_REQUEST)
	) niosv_reset_controller (
		.reset_in0      (reset_in0), // reset_in0.reset
		.reset_in1      (reset_in1), // reset_in1.reset
		.clk            (clk),       //       clk.clk
		.reset_out      (reset_out), // reset_out.reset
		.reset_req      (),          // (terminated)
		.reset_req_in0  (1'b0),      // (terminated)
		.reset_req_in1  (1'b0),      // (terminated)
		.reset_in2      (1'b0),      // (terminated)
		.reset_req_in2  (1'b0),      // (terminated)
		.reset_in3      (1'b0),      // (terminated)
		.reset_req_in3  (1'b0),      // (terminated)
		.reset_in4      (1'b0),      // (terminated)
		.reset_req_in4  (1'b0),      // (terminated)
		.reset_in5      (1'b0),      // (terminated)
		.reset_req_in5  (1'b0),      // (terminated)
		.reset_in6      (1'b0),      // (terminated)
		.reset_req_in6  (1'b0),      // (terminated)
		.reset_in7      (1'b0),      // (terminated)
		.reset_req_in7  (1'b0),      // (terminated)
		.reset_in8      (1'b0),      // (terminated)
		.reset_req_in8  (1'b0),      // (terminated)
		.reset_in9      (1'b0),      // (terminated)
		.reset_req_in9  (1'b0),      // (terminated)
		.reset_in10     (1'b0),      // (terminated)
		.reset_req_in10 (1'b0),      // (terminated)
		.reset_in11     (1'b0),      // (terminated)
		.reset_req_in11 (1'b0),      // (terminated)
		.reset_in12     (1'b0),      // (terminated)
		.reset_req_in12 (1'b0),      // (terminated)
		.reset_in13     (1'b0),      // (terminated)
		.reset_req_in13 (1'b0),      // (terminated)
		.reset_in14     (1'b0),      // (terminated)
		.reset_req_in14 (1'b0),      // (terminated)
		.reset_in15     (1'b0),      // (terminated)
		.reset_req_in15 (1'b0)       // (terminated)
	);

endmodule

// nios.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module nios (
		input  wire       clk_clk,                          //                       clk.clk
		output wire [9:0] pio_0_external_connection_export, // pio_0_external_connection.export
		input  wire       reset_reset_n                     //                     reset.reset_n
	);

	wire  [31:0] intel_niosv_m_0_data_manager_awaddr;                            // intel_niosv_m_0:data_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_awaddr
	wire   [1:0] intel_niosv_m_0_data_manager_bresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_bresp -> intel_niosv_m_0:data_manager_bresp
	wire         intel_niosv_m_0_data_manager_arready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_arready -> intel_niosv_m_0:data_manager_arready
	wire  [31:0] intel_niosv_m_0_data_manager_rdata;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rdata -> intel_niosv_m_0:data_manager_rdata
	wire   [3:0] intel_niosv_m_0_data_manager_wstrb;                             // intel_niosv_m_0:data_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_data_manager_wstrb
	wire         intel_niosv_m_0_data_manager_wready;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_wready -> intel_niosv_m_0:data_manager_wready
	wire         intel_niosv_m_0_data_manager_awready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_awready -> intel_niosv_m_0:data_manager_awready
	wire         intel_niosv_m_0_data_manager_rready;                            // intel_niosv_m_0:data_manager_rready -> mm_interconnect_0:intel_niosv_m_0_data_manager_rready
	wire         intel_niosv_m_0_data_manager_bready;                            // intel_niosv_m_0:data_manager_bready -> mm_interconnect_0:intel_niosv_m_0_data_manager_bready
	wire         intel_niosv_m_0_data_manager_wvalid;                            // intel_niosv_m_0:data_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_wvalid
	wire  [31:0] intel_niosv_m_0_data_manager_araddr;                            // intel_niosv_m_0:data_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_araddr
	wire   [2:0] intel_niosv_m_0_data_manager_arprot;                            // intel_niosv_m_0:data_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_arprot
	wire   [1:0] intel_niosv_m_0_data_manager_rresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rresp -> intel_niosv_m_0:data_manager_rresp
	wire   [2:0] intel_niosv_m_0_data_manager_awprot;                            // intel_niosv_m_0:data_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_awprot
	wire  [31:0] intel_niosv_m_0_data_manager_wdata;                             // intel_niosv_m_0:data_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_data_manager_wdata
	wire         intel_niosv_m_0_data_manager_arvalid;                           // intel_niosv_m_0:data_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_arvalid
	wire         intel_niosv_m_0_data_manager_bvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_bvalid -> intel_niosv_m_0:data_manager_bvalid
	wire         intel_niosv_m_0_data_manager_awvalid;                           // intel_niosv_m_0:data_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_awvalid
	wire         intel_niosv_m_0_data_manager_rvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_rvalid -> intel_niosv_m_0:data_manager_rvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_awaddr;                     // intel_niosv_m_0:instruction_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awaddr
	wire   [1:0] intel_niosv_m_0_instruction_manager_bresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bresp -> intel_niosv_m_0:instruction_manager_bresp
	wire         intel_niosv_m_0_instruction_manager_arready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_arready -> intel_niosv_m_0:instruction_manager_arready
	wire  [31:0] intel_niosv_m_0_instruction_manager_rdata;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rdata -> intel_niosv_m_0:instruction_manager_rdata
	wire   [3:0] intel_niosv_m_0_instruction_manager_wstrb;                      // intel_niosv_m_0:instruction_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wstrb
	wire         intel_niosv_m_0_instruction_manager_wready;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_wready -> intel_niosv_m_0:instruction_manager_wready
	wire         intel_niosv_m_0_instruction_manager_awready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_awready -> intel_niosv_m_0:instruction_manager_awready
	wire         intel_niosv_m_0_instruction_manager_rready;                     // intel_niosv_m_0:instruction_manager_rready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_rready
	wire         intel_niosv_m_0_instruction_manager_bready;                     // intel_niosv_m_0:instruction_manager_bready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_bready
	wire         intel_niosv_m_0_instruction_manager_wvalid;                     // intel_niosv_m_0:instruction_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_araddr;                     // intel_niosv_m_0:instruction_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_araddr
	wire   [2:0] intel_niosv_m_0_instruction_manager_arprot;                     // intel_niosv_m_0:instruction_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arprot
	wire   [1:0] intel_niosv_m_0_instruction_manager_rresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rresp -> intel_niosv_m_0:instruction_manager_rresp
	wire   [2:0] intel_niosv_m_0_instruction_manager_awprot;                     // intel_niosv_m_0:instruction_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awprot
	wire  [31:0] intel_niosv_m_0_instruction_manager_wdata;                      // intel_niosv_m_0:instruction_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wdata
	wire         intel_niosv_m_0_instruction_manager_arvalid;                    // intel_niosv_m_0:instruction_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arvalid
	wire         intel_niosv_m_0_instruction_manager_bvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bvalid -> intel_niosv_m_0:instruction_manager_bvalid
	wire         intel_niosv_m_0_instruction_manager_awvalid;                    // intel_niosv_m_0:instruction_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awvalid
	wire         intel_niosv_m_0_instruction_manager_rvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rvalid -> intel_niosv_m_0:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata;            // intel_niosv_m_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest;         // intel_niosv_m_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_address;             // mm_interconnect_0:intel_niosv_m_0_dm_agent_address -> intel_niosv_m_0:dm_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_read;                // mm_interconnect_0:intel_niosv_m_0_dm_agent_read -> intel_niosv_m_0:dm_agent_read
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid;       // intel_niosv_m_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_write;               // mm_interconnect_0:intel_niosv_m_0_dm_agent_write -> intel_niosv_m_0:dm_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata;           // mm_interconnect_0:intel_niosv_m_0_dm_agent_writedata -> intel_niosv_m_0:dm_agent_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_pio_0_s1_chipselect;                          // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                            // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                             // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                               // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                           // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata;      // intel_niosv_m_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest;   // intel_niosv_m_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address;       // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_address -> intel_niosv_m_0:timer_sw_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read;          // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_read -> intel_niosv_m_0:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable;    // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_byteenable -> intel_niosv_m_0:timer_sw_agent_byteenable
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid; // intel_niosv_m_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write;         // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_write -> intel_niosv_m_0:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata;     // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_writedata -> intel_niosv_m_0:timer_sw_agent_writedata
	wire  [15:0] intel_niosv_m_0_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> intel_niosv_m_0:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [intel_niosv_m_0:ndm_reset_in_reset, intel_niosv_m_0:reset_reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:intel_niosv_m_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, pio_0:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         intel_niosv_m_0_dbg_reset_out_reset;                            // intel_niosv_m_0:dbg_reset_out_reset -> rst_controller:reset_in1

	nios_intel_niosv_m_0 intel_niosv_m_0 (
		.clk                          (clk_clk),                                                        //                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                                 //               reset.reset
		.platform_irq_rx_irq          (intel_niosv_m_0_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.ndm_reset_in_reset           (rst_controller_reset_out_reset),                                 //        ndm_reset_in.reset
		.timer_sw_agent_address       (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //      timer_sw_agent.address
		.timer_sw_agent_byteenable    (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_read          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_write         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                    .write
		.timer_sw_agent_writedata     (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_waitrequest   (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                    .waitrequest
		.timer_sw_agent_readdatavalid (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.instruction_manager_awaddr   (intel_niosv_m_0_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awprot   (intel_niosv_m_0_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (intel_niosv_m_0_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (intel_niosv_m_0_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (intel_niosv_m_0_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (intel_niosv_m_0_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (intel_niosv_m_0_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (intel_niosv_m_0_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (intel_niosv_m_0_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (intel_niosv_m_0_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (intel_niosv_m_0_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (intel_niosv_m_0_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (intel_niosv_m_0_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (intel_niosv_m_0_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (intel_niosv_m_0_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (intel_niosv_m_0_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (intel_niosv_m_0_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (intel_niosv_m_0_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (intel_niosv_m_0_instruction_manager_rready),                     //                    .rready
		.data_manager_awaddr          (intel_niosv_m_0_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awprot          (intel_niosv_m_0_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (intel_niosv_m_0_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (intel_niosv_m_0_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (intel_niosv_m_0_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (intel_niosv_m_0_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (intel_niosv_m_0_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (intel_niosv_m_0_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (intel_niosv_m_0_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (intel_niosv_m_0_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (intel_niosv_m_0_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (intel_niosv_m_0_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (intel_niosv_m_0_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (intel_niosv_m_0_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (intel_niosv_m_0_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (intel_niosv_m_0_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (intel_niosv_m_0_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (intel_niosv_m_0_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (intel_niosv_m_0_data_manager_rready),                            //                    .rready
		.dm_agent_address             (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //            dm_agent.address
		.dm_agent_read                (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                    .readdata
		.dm_agent_write               (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                    .write
		.dm_agent_writedata           (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                    .writedata
		.dm_agent_waitrequest         (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                    .waitrequest
		.dm_agent_readdatavalid       (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //                    .readdatavalid
		.dbg_reset_out_reset          (intel_niosv_m_0_dbg_reset_out_reset)                             //       dbg_reset_out.reset
	);

	altera_avalon_jtag_uart #(
		.readBufferDepth            (64),
		.readIRQThreshold           (8),
		.useRegistersForReadBuffer  (0),
		.useRegistersForWriteBuffer (0),
		.writeBufferDepth           (64),
		.writeIRQThreshold          (8),
		.printingMethod             (0),
		.FIFO_WIDTH                 (8),
		.WR_WIDTHU                  (6),
		.RD_WIDTHU                  (6),
		.write_le                   ("ON"),
		.read_le                    ("ON"),
		.HEX_WRITE_DEPTH_STR        (64),
		.HEX_READ_DEPTH_STR         (64),
		.legacySignalAllow          (0)
	) jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         ()                                                             //               irq.irq
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	nios_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)       // external_connection.export
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.intel_niosv_m_0_data_manager_awaddr               (intel_niosv_m_0_data_manager_awaddr),                            //                intel_niosv_m_0_data_manager.awaddr
		.intel_niosv_m_0_data_manager_awprot               (intel_niosv_m_0_data_manager_awprot),                            //                                            .awprot
		.intel_niosv_m_0_data_manager_awvalid              (intel_niosv_m_0_data_manager_awvalid),                           //                                            .awvalid
		.intel_niosv_m_0_data_manager_awready              (intel_niosv_m_0_data_manager_awready),                           //                                            .awready
		.intel_niosv_m_0_data_manager_wdata                (intel_niosv_m_0_data_manager_wdata),                             //                                            .wdata
		.intel_niosv_m_0_data_manager_wstrb                (intel_niosv_m_0_data_manager_wstrb),                             //                                            .wstrb
		.intel_niosv_m_0_data_manager_wvalid               (intel_niosv_m_0_data_manager_wvalid),                            //                                            .wvalid
		.intel_niosv_m_0_data_manager_wready               (intel_niosv_m_0_data_manager_wready),                            //                                            .wready
		.intel_niosv_m_0_data_manager_bresp                (intel_niosv_m_0_data_manager_bresp),                             //                                            .bresp
		.intel_niosv_m_0_data_manager_bvalid               (intel_niosv_m_0_data_manager_bvalid),                            //                                            .bvalid
		.intel_niosv_m_0_data_manager_bready               (intel_niosv_m_0_data_manager_bready),                            //                                            .bready
		.intel_niosv_m_0_data_manager_araddr               (intel_niosv_m_0_data_manager_araddr),                            //                                            .araddr
		.intel_niosv_m_0_data_manager_arprot               (intel_niosv_m_0_data_manager_arprot),                            //                                            .arprot
		.intel_niosv_m_0_data_manager_arvalid              (intel_niosv_m_0_data_manager_arvalid),                           //                                            .arvalid
		.intel_niosv_m_0_data_manager_arready              (intel_niosv_m_0_data_manager_arready),                           //                                            .arready
		.intel_niosv_m_0_data_manager_rdata                (intel_niosv_m_0_data_manager_rdata),                             //                                            .rdata
		.intel_niosv_m_0_data_manager_rresp                (intel_niosv_m_0_data_manager_rresp),                             //                                            .rresp
		.intel_niosv_m_0_data_manager_rvalid               (intel_niosv_m_0_data_manager_rvalid),                            //                                            .rvalid
		.intel_niosv_m_0_data_manager_rready               (intel_niosv_m_0_data_manager_rready),                            //                                            .rready
		.intel_niosv_m_0_instruction_manager_awaddr        (intel_niosv_m_0_instruction_manager_awaddr),                     //         intel_niosv_m_0_instruction_manager.awaddr
		.intel_niosv_m_0_instruction_manager_awprot        (intel_niosv_m_0_instruction_manager_awprot),                     //                                            .awprot
		.intel_niosv_m_0_instruction_manager_awvalid       (intel_niosv_m_0_instruction_manager_awvalid),                    //                                            .awvalid
		.intel_niosv_m_0_instruction_manager_awready       (intel_niosv_m_0_instruction_manager_awready),                    //                                            .awready
		.intel_niosv_m_0_instruction_manager_wdata         (intel_niosv_m_0_instruction_manager_wdata),                      //                                            .wdata
		.intel_niosv_m_0_instruction_manager_wstrb         (intel_niosv_m_0_instruction_manager_wstrb),                      //                                            .wstrb
		.intel_niosv_m_0_instruction_manager_wvalid        (intel_niosv_m_0_instruction_manager_wvalid),                     //                                            .wvalid
		.intel_niosv_m_0_instruction_manager_wready        (intel_niosv_m_0_instruction_manager_wready),                     //                                            .wready
		.intel_niosv_m_0_instruction_manager_bresp         (intel_niosv_m_0_instruction_manager_bresp),                      //                                            .bresp
		.intel_niosv_m_0_instruction_manager_bvalid        (intel_niosv_m_0_instruction_manager_bvalid),                     //                                            .bvalid
		.intel_niosv_m_0_instruction_manager_bready        (intel_niosv_m_0_instruction_manager_bready),                     //                                            .bready
		.intel_niosv_m_0_instruction_manager_araddr        (intel_niosv_m_0_instruction_manager_araddr),                     //                                            .araddr
		.intel_niosv_m_0_instruction_manager_arprot        (intel_niosv_m_0_instruction_manager_arprot),                     //                                            .arprot
		.intel_niosv_m_0_instruction_manager_arvalid       (intel_niosv_m_0_instruction_manager_arvalid),                    //                                            .arvalid
		.intel_niosv_m_0_instruction_manager_arready       (intel_niosv_m_0_instruction_manager_arready),                    //                                            .arready
		.intel_niosv_m_0_instruction_manager_rdata         (intel_niosv_m_0_instruction_manager_rdata),                      //                                            .rdata
		.intel_niosv_m_0_instruction_manager_rresp         (intel_niosv_m_0_instruction_manager_rresp),                      //                                            .rresp
		.intel_niosv_m_0_instruction_manager_rvalid        (intel_niosv_m_0_instruction_manager_rvalid),                     //                                            .rvalid
		.intel_niosv_m_0_instruction_manager_rready        (intel_niosv_m_0_instruction_manager_rready),                     //                                            .rready
		.clk_0_clk_clk                                     (clk_clk),                                                        //                                   clk_0_clk.clk
		.intel_niosv_m_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // intel_niosv_m_0_reset_reset_bridge_in_reset.reset
		.intel_niosv_m_0_dm_agent_address                  (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //                    intel_niosv_m_0_dm_agent.address
		.intel_niosv_m_0_dm_agent_write                    (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                                            .write
		.intel_niosv_m_0_dm_agent_read                     (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                                            .read
		.intel_niosv_m_0_dm_agent_readdata                 (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                                            .readdata
		.intel_niosv_m_0_dm_agent_writedata                (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                                            .writedata
		.intel_niosv_m_0_dm_agent_readdatavalid            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //                                            .readdatavalid
		.intel_niosv_m_0_dm_agent_waitrequest              (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                                            .waitrequest
		.intel_niosv_m_0_timer_sw_agent_address            (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //              intel_niosv_m_0_timer_sw_agent.address
		.intel_niosv_m_0_timer_sw_agent_write              (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                                            .write
		.intel_niosv_m_0_timer_sw_agent_read               (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                                            .read
		.intel_niosv_m_0_timer_sw_agent_readdata           (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                                            .readdata
		.intel_niosv_m_0_timer_sw_agent_writedata          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                                            .writedata
		.intel_niosv_m_0_timer_sw_agent_byteenable         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                                            .byteenable
		.intel_niosv_m_0_timer_sw_agent_readdatavalid      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                                            .readdatavalid
		.intel_niosv_m_0_timer_sw_agent_waitrequest        (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                            .chipselect
		.onchip_memory2_0_s1_address                       (mm_interconnect_0_onchip_memory2_0_s1_address),                  //                         onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                         (mm_interconnect_0_onchip_memory2_0_s1_write),                    //                                            .write
		.onchip_memory2_0_s1_readdata                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                 //                                            .readdata
		.onchip_memory2_0_s1_writedata                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                //                                            .writedata
		.onchip_memory2_0_s1_byteenable                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),               //                                            .byteenable
		.onchip_memory2_0_s1_chipselect                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),               //                                            .chipselect
		.onchip_memory2_0_s1_clken                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                    //                                            .clken
		.pio_0_s1_address                                  (mm_interconnect_0_pio_0_s1_address),                             //                                    pio_0_s1.address
		.pio_0_s1_write                                    (mm_interconnect_0_pio_0_s1_write),                               //                                            .write
		.pio_0_s1_readdata                                 (mm_interconnect_0_pio_0_s1_readdata),                            //                                            .readdata
		.pio_0_s1_writedata                                (mm_interconnect_0_pio_0_s1_writedata),                           //                                            .writedata
		.pio_0_s1_chipselect                               (mm_interconnect_0_pio_0_s1_chipselect)                           //                                            .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk        (clk_clk),                             //       clk.clk
		.reset      (rst_controller_reset_out_reset),      // clk_reset.reset
		.sender_irq (intel_niosv_m_0_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (intel_niosv_m_0_dbg_reset_out_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
